`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "ahb_cfg.sv"
`include "ahb_slave.sv"
`include "ahb_intf.sv"
`include "ahb_tx.sv"
`include "ahb_seq.sv"
`include "ahb_sqr.sv"
`include "ahb_dvr.sv"
`include "ahb_mon.sv"
`include "ahb_cov.sv"
`include "ahb_master_agent.sv"
//`include "ahb_slave.sv"
`include "ahb_env.sv"
`include "ahb_top.sv"
