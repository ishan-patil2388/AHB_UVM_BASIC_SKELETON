
class ahb_sqr extends uvm_sequencer#(ahb_tx);
	`uvm_component_utils(ahb_sqr)
	`NEW_COMP

		
endclass :ahb_sqr
